module adder(A, B, CI, Y, C, V);

  // inputs
  input [7:0] A, B;
  input CI;

  // outputs
  output [7:0] Y;
  output C, V;

  /* ADD YOUR CODE BELOW THIS LINE */

  /* ADD YOUR CODE ABOVE THIS LINE */


endmodule
